interface SPI_Wrapper_GM_if();

logic MISO_gm;
endinterface