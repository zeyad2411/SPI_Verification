module ;