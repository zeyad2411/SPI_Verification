package shared_pkg;

typedef enum bit [1:0] { WA = 2'b00 , WD = 2'b01 , RA = 2'b10 , RD = 2'b11  } rw_e;
endpackage